*

.SUBCKT		Cadence_Demo_091724_163748_8672
+			J5_1
+			J5_4
+			J6_A1
+			J6_A23
+			J6_C1
+			J6_D3
+			J7_137
+			J7_99
+			LCD1_1
+			LCD1_2
+			LCD2_1
+			LCD2_2
+			P1_1
+			P1_12
+			P1_14
+			P1_2
+			P1_4
+			P1_6
+			U10_11
+			U10_18
+			U10_20
+			U11_11
+			U11_18
+			U11_20
+			U12_A9
+			U12_J2
+			U12_N1
+			U13_A1
+			U13_B2
+			U13_J2
+			U1_D15
+			U1_K10
+			U1_R4
+			U1_T1
+			U22_1
+			U22_20
+			U29_A1
+			U29_H5
+			U29_J1
+			U29_L7
+			U2_A16
+			U2_B13
+			U2_K10
+			U2_K13
+			U2_R8
+			U30_A1
+			U30_A5
+			U30_H5
+			U30_J1
+			U31_A1
+			U31_J1
+			U31_L7
+			U32_10
+			U32_2
+			U33_3
+			U33_4
+			U33_7
+			U35_10
+			U35_9
+			U36_3
+			U36_4
+			U36_7
+			U38_1
+			U38_20
+			U39_1
+			U39_20
+			U3_3
+			U3_8
+			U40_16
+			U40_32
+			U41_16
+			U41_32
+			U42_24
+			U42_32
+			U43_24
+			U43_32
+			U44_24
+			U44_32
+			U45_16
+			U45_32
+			U46_16
+			U46_32
+			U47_16
+			U47_32
+			U48_10
+			U48_20
+			U49_1
+			U49_4
+			U50_1
+			U50_28
+			U51_10
+			U51_2
+			U51_5
+			U51_8
+			U5_1
+			U5_4
+			U6_25
+			U6_42
+			U7_10
+			U7_20
+			U8_34
+			U8_42
+			U9_4
+			U9_42
*The following is the Cadence MCP(model connection protocol) Section
***********************************
*[MCP Begin]
*[MCP Ver] 1.2
*[MCP Source] Cadence Design Systems, Inc. MCP Editor
*
*[REM]***********************************************************************
*[Connection] J5 USB3A_FEMALE_USB3A_FEMALE_IO_AU-Y1005-3-R_PSL-00000013_AU-Y1005-3-R 3
*[Connection Type] 
*[Power Nets]
*1	J5_1	VCC	0.095550000000	0.057300000000
*[Ground Nets]
*4	J5_4	GND_DIGITAL	0.095550000000	0.064300000000
*7	J5_4	GND_DIGITAL	0.094050000000	0.060800000000
*
*
*[REM]***********************************************************************
*[Connection] J6 CONN_C1367550_6_C-1367550-6_IO_(S1+S2+S3+S4+S5+S6)_6367550-6_PSL-00000038_6367550-6 20
*[Connection Type] 
*[Power Nets]
*A1	J6_A1	V+12	-0.012784000000	0.023255000000
*A2	J6_A1	V+12	-0.012784000000	0.025285000000
*D1	J6_A1	V+12	-0.018784000000	0.023255000000
*D2	J6_A1	V+12	-0.018784000000	0.025285000000
*A23	J6_A23	VCC	-0.012784000000	0.079135000000
*A24	J6_A23	VCC	-0.012784000000	0.081165000000
*D23	J6_A23	VCC	-0.018784000000	0.079135000000
*D24	J6_A23	VCC	-0.018784000000	0.081165000000
*A3	J6_D3	V12N	-0.012784000000	0.028335000000
*A4	J6_D3	V12N	-0.012784000000	0.030365000000
*D3	J6_D3	V12N	-0.018784000000	0.028335000000
*D4	J6_D3	V12N	-0.018784000000	0.030365000000
*[Ground Nets]
*C1	J6_C1	GND_DIGITAL	-0.016284000000	0.025795000000
*C2	J6_C1	GND_DIGITAL	-0.016284000000	0.027825000000
*C23	J6_C1	GND_DIGITAL	-0.016284000000	0.081675000000
*C24	J6_C1	GND_DIGITAL	-0.016284000000	0.083705000000
*F1	J6_C1	GND_DIGITAL	-0.022284000000	0.025795000000
*F2	J6_C1	GND_DIGITAL	-0.022284000000	0.027825000000
*F23	J6_C1	GND_DIGITAL	-0.022284000000	0.081675000000
*F24	J6_C1	GND_DIGITAL	-0.022284000000	0.083705000000
*
*
*[REM]***********************************************************************
*[Connection] J7 CONN_DIMM_200_C_1_1473005_1_J1_IO_(S1+S2+S3+S4)_1473005-1_PSL-00000043_1473005-1 80
*[Connection Type] 
*[Power Nets]
*131	J7_137	VCC	0.052550000000	0.101650000000
*132	J7_137	VCC	0.052850000000	0.093450000000
*133	J7_137	VCC	0.053150000000	0.101650000000
*134	J7_137	VCC	0.053450000000	0.093450000000
*135	J7_137	VCC	0.053750000000	0.101650000000
*136	J7_137	VCC	0.054050000000	0.093450000000
*137	J7_137	VCC	0.054350000000	0.101650000000
*138	J7_137	VCC	0.054650000000	0.093450000000
*181	J7_137	VCC	0.067550000000	0.101650000000
*182	J7_137	VCC	0.067850000000	0.093450000000
*183	J7_137	VCC	0.068150000000	0.101650000000
*184	J7_137	VCC	0.068450000000	0.093450000000
*185	J7_137	VCC	0.068750000000	0.101650000000
*186	J7_137	VCC	0.069050000000	0.093450000000
*187	J7_137	VCC	0.069350000000	0.101650000000
*188	J7_137	VCC	0.069650000000	0.093450000000
*31	J7_137	VCC	0.018950000000	0.101650000000
*32	J7_137	VCC	0.019250000000	0.093450000000
*33	J7_137	VCC	0.019550000000	0.101650000000
*34	J7_137	VCC	0.019850000000	0.093450000000
*35	J7_137	VCC	0.020150000000	0.101650000000
*36	J7_137	VCC	0.020450000000	0.093450000000
*37	J7_137	VCC	0.020750000000	0.101650000000
*38	J7_137	VCC	0.021050000000	0.093450000000
*81	J7_137	VCC	0.037550000000	0.101650000000
*82	J7_137	VCC	0.037850000000	0.093450000000
*83	J7_137	VCC	0.038150000000	0.101650000000
*84	J7_137	VCC	0.038450000000	0.093450000000
*85	J7_137	VCC	0.038750000000	0.101650000000
*86	J7_137	VCC	0.039050000000	0.093450000000
*87	J7_137	VCC	0.039350000000	0.101650000000
*88	J7_137	VCC	0.039650000000	0.093450000000
*[Ground Nets]
*100	J7_99	GND_DIGITAL	0.043250000000	0.093450000000
*139	J7_99	GND_DIGITAL	0.054950000000	0.101650000000
*140	J7_99	GND_DIGITAL	0.055250000000	0.093450000000
*141	J7_99	GND_DIGITAL	0.055550000000	0.101650000000
*142	J7_99	GND_DIGITAL	0.055850000000	0.093450000000
*143	J7_99	GND_DIGITAL	0.056150000000	0.101650000000
*144	J7_99	GND_DIGITAL	0.056450000000	0.093450000000
*145	J7_99	GND_DIGITAL	0.056750000000	0.101650000000
*146	J7_99	GND_DIGITAL	0.057050000000	0.093450000000
*147	J7_99	GND_DIGITAL	0.057350000000	0.101650000000
*148	J7_99	GND_DIGITAL	0.057650000000	0.093450000000
*149	J7_99	GND_DIGITAL	0.057950000000	0.101650000000
*150	J7_99	GND_DIGITAL	0.058250000000	0.093450000000
*189	J7_99	GND_DIGITAL	0.069950000000	0.101650000000
*190	J7_99	GND_DIGITAL	0.070250000000	0.093450000000
*191	J7_99	GND_DIGITAL	0.070550000000	0.101650000000
*192	J7_99	GND_DIGITAL	0.070850000000	0.093450000000
*193	J7_99	GND_DIGITAL	0.071150000000	0.101650000000
*194	J7_99	GND_DIGITAL	0.071450000000	0.093450000000
*195	J7_99	GND_DIGITAL	0.071750000000	0.101650000000
*196	J7_99	GND_DIGITAL	0.072050000000	0.093450000000
*197	J7_99	GND_DIGITAL	0.072350000000	0.101650000000
*198	J7_99	GND_DIGITAL	0.072650000000	0.093450000000
*199	J7_99	GND_DIGITAL	0.072950000000	0.101650000000
*200	J7_99	GND_DIGITAL	0.073250000000	0.093450000000
*39	J7_99	GND_DIGITAL	0.021350000000	0.101650000000
*40	J7_99	GND_DIGITAL	0.021650000000	0.093450000000
*41	J7_99	GND_DIGITAL	0.025550000000	0.101650000000
*42	J7_99	GND_DIGITAL	0.025850000000	0.093450000000
*43	J7_99	GND_DIGITAL	0.026150000000	0.101650000000
*44	J7_99	GND_DIGITAL	0.026450000000	0.093450000000
*45	J7_99	GND_DIGITAL	0.026750000000	0.101650000000
*46	J7_99	GND_DIGITAL	0.027050000000	0.093450000000
*47	J7_99	GND_DIGITAL	0.027350000000	0.101650000000
*48	J7_99	GND_DIGITAL	0.027650000000	0.093450000000
*49	J7_99	GND_DIGITAL	0.027950000000	0.101650000000
*50	J7_99	GND_DIGITAL	0.028250000000	0.093450000000
*89	J7_99	GND_DIGITAL	0.039950000000	0.101650000000
*90	J7_99	GND_DIGITAL	0.040250000000	0.093450000000
*91	J7_99	GND_DIGITAL	0.040550000000	0.101650000000
*92	J7_99	GND_DIGITAL	0.040850000000	0.093450000000
*93	J7_99	GND_DIGITAL	0.041150000000	0.101650000000
*94	J7_99	GND_DIGITAL	0.041450000000	0.093450000000
*95	J7_99	GND_DIGITAL	0.041750000000	0.101650000000
*96	J7_99	GND_DIGITAL	0.042050000000	0.093450000000
*97	J7_99	GND_DIGITAL	0.042350000000	0.101650000000
*98	J7_99	GND_DIGITAL	0.042650000000	0.093450000000
*99	J7_99	GND_DIGITAL	0.042950000000	0.101650000000
*
*
*[REM]***********************************************************************
*[Connection] LCD1 LCD-EA-8081-A3N_LCD_EA_8081-A3N-B_DISCRETE_S1D13742F01A200_PSL-00000046_S1D13742F01A200 3
*[Connection Type] 
*[Power Nets]
*2	LCD1_2	VCC	0.026200000000	0.173060000000
*[Ground Nets]
*1	LCD1_1	GND_DIGITAL	0.026200000000	0.175600000000
*3	LCD1_1	GND_DIGITAL	0.026200000000	0.170520000000
*
*
*[REM]***********************************************************************
*[Connection] LCD2 LCD-EA-8081-A3N_LCD_EA_8081-A3N-B_DISCRETE_S1D13742F01A200_PSL-00000046_S1D13742F01A200 3
*[Connection Type] 
*[Power Nets]
*2	LCD2_2	VCC	0.067700000000	0.173060000000
*[Ground Nets]
*1	LCD2_1	GND_DIGITAL	0.067700000000	0.175600000000
*3	LCD2_1	GND_DIGITAL	0.067700000000	0.170520000000
*
*
*[REM]***********************************************************************
*[Connection] P1 HDR_2X7_M_SAMTEC_TST-107-XX-X-D_IO_TST-107-01-G-D_EMA-00006288V22_TST-107-01-G-D 9
*[Connection Type] 
*[Power Nets]
*12	P1_12	3V3	0.012200000000	0.025860000000
*14	P1_14	2V5	0.009660000000	0.025860000000
*2	P1_2	0V9	0.024900000000	0.025860000000
*4	P1_4	1V2	0.022360000000	0.025860000000
*6	P1_6	1V8	0.019820000000	0.025860000000
*[Ground Nets]
*1	P1_1	GND_DIGITAL	0.024900000000	0.028400000000
*13	P1_1	GND_DIGITAL	0.009660000000	0.028400000000
*5	P1_1	GND_DIGITAL	0.019820000000	0.028400000000
*9	P1_1	GND_DIGITAL	0.014740000000	0.028400000000
*
*
*[REM]***********************************************************************
*[Connection] U1 DEMOG_INTERFACE_FT256_IC_(S1+S2+S3+S4+S5+S6)_XC6SLX25-3FTG256_PSL-00000032_XC6SLX25-3FTG256 62
*[Connection Type] 
*[Power Nets]
*B13	U1_D15	3V3	0.017000000000	0.068000000000
*B4	U1_D15	3V3	0.026000000000	0.068000000000
*B9	U1_D15	3V3	0.021000000000	0.068000000000
*D10	U1_D15	3V3	0.020000000000	0.070000000000
*D15	U1_D15	3V3	0.015000000000	0.070000000000
*D7	U1_D15	3V3	0.023000000000	0.070000000000
*G13	U1_D15	3V3	0.017000000000	0.073000000000
*J15	U1_D15	3V3	0.015000000000	0.075000000000
*K13	U1_D15	3V3	0.017000000000	0.076000000000
*N15	U1_D15	3V3	0.015000000000	0.079000000000
*G7	U1_K10	1V2	0.023000000000	0.073000000000
*G9	U1_K10	1V2	0.021000000000	0.073000000000
*H10	U1_K10	1V2	0.020000000000	0.074000000000
*H8	U1_K10	1V2	0.022000000000	0.074000000000
*J7	U1_K10	1V2	0.023000000000	0.075000000000
*J9	U1_K10	1V2	0.021000000000	0.075000000000
*K10	U1_K10	1V2	0.020000000000	0.076000000000
*K8	U1_K10	1V2	0.022000000000	0.076000000000
*D2	U1_R4	2V5	0.028000000000	0.070000000000
*E5	U1_R4	2V5	0.025000000000	0.071000000000
*F11	U1_R4	2V5	0.019000000000	0.072000000000
*F8	U1_R4	2V5	0.022000000000	0.072000000000
*G10	U1_R4	2V5	0.020000000000	0.073000000000
*G4	U1_R4	2V5	0.026000000000	0.073000000000
*H6	U1_R4	2V5	0.024000000000	0.074000000000
*J10	U1_R4	2V5	0.020000000000	0.075000000000
*J2	U1_R4	2V5	0.028000000000	0.075000000000
*K4	U1_R4	2V5	0.026000000000	0.076000000000
*L6	U1_R4	2V5	0.024000000000	0.077000000000
*L9	U1_R4	2V5	0.021000000000	0.077000000000
*N10	U1_R4	2V5	0.020000000000	0.079000000000
*N2	U1_R4	2V5	0.028000000000	0.079000000000
*N7	U1_R4	2V5	0.023000000000	0.079000000000
*R13	U1_R4	2V5	0.017000000000	0.081000000000
*R4	U1_R4	2V5	0.026000000000	0.081000000000
*R8	U1_R4	2V5	0.022000000000	0.081000000000
*[Ground Nets]
*A1	U1_T1	GND_DIGITAL	0.029000000000	0.067000000000
*A16	U1_T1	GND_DIGITAL	0.014000000000	0.067000000000
*B11	U1_T1	GND_DIGITAL	0.019000000000	0.068000000000
*B7	U1_T1	GND_DIGITAL	0.023000000000	0.068000000000
*D13	U1_T1	GND_DIGITAL	0.017000000000	0.070000000000
*D4	U1_T1	GND_DIGITAL	0.026000000000	0.070000000000
*E9	U1_T1	GND_DIGITAL	0.021000000000	0.071000000000
*G15	U1_T1	GND_DIGITAL	0.015000000000	0.073000000000
*G2	U1_T1	GND_DIGITAL	0.028000000000	0.073000000000
*G8	U1_T1	GND_DIGITAL	0.022000000000	0.073000000000
*H12	U1_T1	GND_DIGITAL	0.018000000000	0.074000000000
*H7	U1_T1	GND_DIGITAL	0.023000000000	0.074000000000
*H9	U1_T1	GND_DIGITAL	0.021000000000	0.074000000000
*J5	U1_T1	GND_DIGITAL	0.025000000000	0.075000000000
*J8	U1_T1	GND_DIGITAL	0.022000000000	0.075000000000
*K7	U1_T1	GND_DIGITAL	0.023000000000	0.076000000000
*K9	U1_T1	GND_DIGITAL	0.021000000000	0.076000000000
*L15	U1_T1	GND_DIGITAL	0.015000000000	0.077000000000
*L2	U1_T1	GND_DIGITAL	0.028000000000	0.077000000000
*M8	U1_T1	GND_DIGITAL	0.022000000000	0.078000000000
*N13	U1_T1	GND_DIGITAL	0.017000000000	0.079000000000
*P3	U1_T1	GND_DIGITAL	0.027000000000	0.080000000000
*R10	U1_T1	GND_DIGITAL	0.020000000000	0.081000000000
*R6	U1_T1	GND_DIGITAL	0.024000000000	0.081000000000
*T1	U1_T1	GND_DIGITAL	0.029000000000	0.082000000000
*T16	U1_T1	GND_DIGITAL	0.014000000000	0.082000000000
*
*
*[REM]***********************************************************************
*[Connection] U10 XCF01SVOG20_XCF01SVOG20_IC_XCF01SVOG20C_PSL-00000005_XCF01SVOG20C 4
*[Connection Type] 
*[Power Nets]
*18	U10_18	3V3	0.043286000000	0.066903000000
*19	U10_20	2V5	0.043286000000	0.067553000000
*20	U10_20	2V5	0.043286000000	0.068203000000
*[Ground Nets]
*11	U10_11	GND_DIGITAL	0.043286000000	0.062353000000
*
*
*[REM]***********************************************************************
*[Connection] U11 XCF01SVOG20_XCF01SVOG20_IC_XCF01SVOG20C_PSL-00000030_XCF01SVOG20C 4
*[Connection Type] 
*[Power Nets]
*18	U11_18	3V3	0.049400000000	0.045625000000
*19	U11_20	2V5	0.049400000000	0.044975000000
*20	U11_20	2V5	0.049400000000	0.044325000000
*[Ground Nets]
*11	U11_11	GND_DIGITAL	0.049400000000	0.050175000000
*
*
*[REM]***********************************************************************
*[Connection] U12 MT47H64M16_MT47H128M_IC_(S1+S2)_MT47H64M16HR-3:G_TR_PSL-00000002_MT47H64M16HR-3:G_TR 32
*[Connection Type] 
*[Power Nets]
*A1	U12_A9	1V8	0.018100000000	0.056600000000
*A9	U12_A9	1V8	0.018100000000	0.050200000000
*C1	U12_A9	1V8	0.016500000000	0.056600000000
*C3	U12_A9	1V8	0.016500000000	0.055000000000
*C7	U12_A9	1V8	0.016500000000	0.051800000000
*C9	U12_A9	1V8	0.016500000000	0.050200000000
*E1	U12_A9	1V8	0.014900000000	0.056600000000
*E9	U12_A9	1V8	0.014900000000	0.050200000000
*G1	U12_A9	1V8	0.013300000000	0.056600000000
*G7	U12_A9	1V8	0.013300000000	0.051800000000
*G9	U12_A9	1V8	0.013300000000	0.050200000000
*J1	U12_A9	1V8	0.011700000000	0.056600000000
*J9	U12_A9	1V8	0.011700000000	0.050200000000
*M9	U12_A9	1V8	0.009300000000	0.050200000000
*R1	U12_A9	1V8	0.006900000000	0.056600000000
*J2	U12_J2	0V9	0.011700000000	0.055800000000
*[Ground Nets]
*A3	U12_N1	GND_DIGITAL	0.018100000000	0.055000000000
*A7	U12_N1	GND_DIGITAL	0.018100000000	0.051800000000
*B2	U12_N1	GND_DIGITAL	0.017300000000	0.055800000000
*B8	U12_N1	GND_DIGITAL	0.017300000000	0.051000000000
*D2	U12_N1	GND_DIGITAL	0.015700000000	0.055800000000
*D8	U12_N1	GND_DIGITAL	0.015700000000	0.051000000000
*E3	U12_N1	GND_DIGITAL	0.014900000000	0.055000000000
*E7	U12_N1	GND_DIGITAL	0.014900000000	0.051800000000
*F2	U12_N1	GND_DIGITAL	0.014100000000	0.055800000000
*F8	U12_N1	GND_DIGITAL	0.014100000000	0.051000000000
*H2	U12_N1	GND_DIGITAL	0.012500000000	0.055800000000
*H8	U12_N1	GND_DIGITAL	0.012500000000	0.051000000000
*J3	U12_N1	GND_DIGITAL	0.011700000000	0.055000000000
*J7	U12_N1	GND_DIGITAL	0.011700000000	0.051800000000
*N1	U12_N1	GND_DIGITAL	0.008500000000	0.056600000000
*P9	U12_N1	GND_DIGITAL	0.007700000000	0.050200000000
*
*
*[REM]***********************************************************************
*[Connection] U13 MT47H64M16_MT47H128M_IC_(S1+S2)_MT47H64M16HR-3:G_TR_PSL-00000002_MT47H64M16HR-3:G_TR 32
*[Connection Type] 
*[Power Nets]
*A1	U13_A1	1V8	0.018100000000	0.042800000000
*A9	U13_A1	1V8	0.018100000000	0.036400000000
*C1	U13_A1	1V8	0.016500000000	0.042800000000
*C3	U13_A1	1V8	0.016500000000	0.041200000000
*C7	U13_A1	1V8	0.016500000000	0.038000000000
*C9	U13_A1	1V8	0.016500000000	0.036400000000
*E1	U13_A1	1V8	0.014900000000	0.042800000000
*E9	U13_A1	1V8	0.014900000000	0.036400000000
*G1	U13_A1	1V8	0.013300000000	0.042800000000
*G7	U13_A1	1V8	0.013300000000	0.038000000000
*G9	U13_A1	1V8	0.013300000000	0.036400000000
*J1	U13_A1	1V8	0.011700000000	0.042800000000
*J9	U13_A1	1V8	0.011700000000	0.036400000000
*M9	U13_A1	1V8	0.009300000000	0.036400000000
*R1	U13_A1	1V8	0.006900000000	0.042800000000
*J2	U13_J2	0V9	0.011700000000	0.042000000000
*[Ground Nets]
*A3	U13_B2	GND_DIGITAL	0.018100000000	0.041200000000
*A7	U13_B2	GND_DIGITAL	0.018100000000	0.038000000000
*B2	U13_B2	GND_DIGITAL	0.017300000000	0.042000000000
*B8	U13_B2	GND_DIGITAL	0.017300000000	0.037200000000
*D2	U13_B2	GND_DIGITAL	0.015700000000	0.042000000000
*D8	U13_B2	GND_DIGITAL	0.015700000000	0.037200000000
*E3	U13_B2	GND_DIGITAL	0.014900000000	0.041200000000
*E7	U13_B2	GND_DIGITAL	0.014900000000	0.038000000000
*F2	U13_B2	GND_DIGITAL	0.014100000000	0.042000000000
*F8	U13_B2	GND_DIGITAL	0.014100000000	0.037200000000
*H2	U13_B2	GND_DIGITAL	0.012500000000	0.042000000000
*H8	U13_B2	GND_DIGITAL	0.012500000000	0.037200000000
*J3	U13_B2	GND_DIGITAL	0.011700000000	0.041200000000
*J7	U13_B2	GND_DIGITAL	0.011700000000	0.038000000000
*N1	U13_B2	GND_DIGITAL	0.008500000000	0.042800000000
*P9	U13_B2	GND_DIGITAL	0.007700000000	0.036400000000
*
*
*[REM]***********************************************************************
*[Connection] U2 DEMOG_COPROC_FT256_IC_(S1+S2+S3+S4+S5+S6)_XC6SLX25-3FTG256_PSL-00000033_XC6SLX25-3FTG256 62
*[Connection Type] 
*[Power Nets]
*B13	U2_B13	1V8	0.038350000000	0.049950000000
*B4	U2_B13	1V8	0.029350000000	0.049950000000
*B9	U2_B13	1V8	0.034350000000	0.049950000000
*D2	U2_B13	1V8	0.027350000000	0.047950000000
*G4	U2_B13	1V8	0.029350000000	0.044950000000
*J2	U2_B13	1V8	0.027350000000	0.042950000000
*K4	U2_B13	1V8	0.029350000000	0.041950000000
*N15	U2_B13	1V8	0.040350000000	0.038950000000
*N2	U2_B13	1V8	0.027350000000	0.038950000000
*N7	U2_B13	1V8	0.032350000000	0.038950000000
*R13	U2_B13	1V8	0.038350000000	0.036950000000
*G7	U2_K10	1V2	0.032350000000	0.044950000000
*G9	U2_K10	1V2	0.034350000000	0.044950000000
*H10	U2_K10	1V2	0.035350000000	0.043950000000
*H8	U2_K10	1V2	0.033350000000	0.043950000000
*J7	U2_K10	1V2	0.032350000000	0.042950000000
*J9	U2_K10	1V2	0.034350000000	0.042950000000
*K10	U2_K10	1V2	0.035350000000	0.041950000000
*K8	U2_K10	1V2	0.033350000000	0.041950000000
*G13	U2_K13	3V3	0.038350000000	0.044950000000
*J15	U2_K13	3V3	0.040350000000	0.042950000000
*K13	U2_K13	3V3	0.038350000000	0.041950000000
*D10	U2_R8	2V5	0.035350000000	0.047950000000
*D15	U2_R8	2V5	0.040350000000	0.047950000000
*D7	U2_R8	2V5	0.032350000000	0.047950000000
*E5	U2_R8	2V5	0.030350000000	0.046950000000
*F11	U2_R8	2V5	0.036350000000	0.045950000000
*F8	U2_R8	2V5	0.033350000000	0.045950000000
*G10	U2_R8	2V5	0.035350000000	0.044950000000
*H6	U2_R8	2V5	0.031350000000	0.043950000000
*J10	U2_R8	2V5	0.035350000000	0.042950000000
*L6	U2_R8	2V5	0.031350000000	0.040950000000
*L9	U2_R8	2V5	0.034350000000	0.040950000000
*N10	U2_R8	2V5	0.035350000000	0.038950000000
*R4	U2_R8	2V5	0.029350000000	0.036950000000
*R8	U2_R8	2V5	0.033350000000	0.036950000000
*[Ground Nets]
*A1	U2_A16	GND_DIGITAL	0.026350000000	0.050950000000
*A16	U2_A16	GND_DIGITAL	0.041350000000	0.050950000000
*B11	U2_A16	GND_DIGITAL	0.036350000000	0.049950000000
*B7	U2_A16	GND_DIGITAL	0.032350000000	0.049950000000
*D13	U2_A16	GND_DIGITAL	0.038350000000	0.047950000000
*D4	U2_A16	GND_DIGITAL	0.029350000000	0.047950000000
*E9	U2_A16	GND_DIGITAL	0.034350000000	0.046950000000
*G15	U2_A16	GND_DIGITAL	0.040350000000	0.044950000000
*G2	U2_A16	GND_DIGITAL	0.027350000000	0.044950000000
*G8	U2_A16	GND_DIGITAL	0.033350000000	0.044950000000
*H12	U2_A16	GND_DIGITAL	0.037350000000	0.043950000000
*H7	U2_A16	GND_DIGITAL	0.032350000000	0.043950000000
*H9	U2_A16	GND_DIGITAL	0.034350000000	0.043950000000
*J5	U2_A16	GND_DIGITAL	0.030350000000	0.042950000000
*J8	U2_A16	GND_DIGITAL	0.033350000000	0.042950000000
*K7	U2_A16	GND_DIGITAL	0.032350000000	0.041950000000
*K9	U2_A16	GND_DIGITAL	0.034350000000	0.041950000000
*L15	U2_A16	GND_DIGITAL	0.040350000000	0.040950000000
*L2	U2_A16	GND_DIGITAL	0.027350000000	0.040950000000
*M8	U2_A16	GND_DIGITAL	0.033350000000	0.039950000000
*N13	U2_A16	GND_DIGITAL	0.038350000000	0.038950000000
*P3	U2_A16	GND_DIGITAL	0.028350000000	0.037950000000
*R10	U2_A16	GND_DIGITAL	0.035350000000	0.036950000000
*R6	U2_A16	GND_DIGITAL	0.031350000000	0.036950000000
*T1	U2_A16	GND_DIGITAL	0.026350000000	0.035950000000
*T16	U2_A16	GND_DIGITAL	0.041350000000	0.035950000000
*
*
*[REM]***********************************************************************
*[Connection] U22 FF_D_8X_OE3S_20P_SOIC127P1032X265-20AN_IC_74HCT574_EMA-00007307V22_74HCT574 3
*[Connection Type] 
*[Power Nets]
*20	U22_20	VCC	0.084250000000	0.041115000000
*[Ground Nets]
*1	U22_1	GND_DIGITAL	0.074750000000	0.041115000000
*10	U22_1	GND_DIGITAL	0.074750000000	0.029685000000
*
*
*[REM]***********************************************************************
*[Connection] U29 LTM8025_LTUMODULE7X11_IC_LTM8025EV#PBF_PSL-00000026_LTM8025EV#PBF 65
*[Connection Type] 
*[Power Nets]
*A1	U29_A1	1V2	0.059436000000	0.059182000000
*A2	U29_A1	1V2	0.060706000000	0.059182000000
*A3	U29_A1	1V2	0.061976000000	0.059182000000
*A4	U29_A1	1V2	0.063246000000	0.059182000000
*B1	U29_A1	1V2	0.059436000000	0.057912000000
*B2	U29_A1	1V2	0.060706000000	0.057912000000
*B3	U29_A1	1V2	0.061976000000	0.057912000000
*B4	U29_A1	1V2	0.063246000000	0.057912000000
*C1	U29_A1	1V2	0.059436000000	0.056642000000
*C2	U29_A1	1V2	0.060706000000	0.056642000000
*C3	U29_A1	1V2	0.061976000000	0.056642000000
*C4	U29_A1	1V2	0.063246000000	0.056642000000
*D1	U29_A1	1V2	0.059436000000	0.055372000000
*D2	U29_A1	1V2	0.060706000000	0.055372000000
*D3	U29_A1	1V2	0.061976000000	0.055372000000
*D4	U29_A1	1V2	0.063246000000	0.055372000000
*H5	U29_H5	3V3	0.064516000000	0.050292000000
*J1	U29_J1	V+12	0.059436000000	0.049022000000
*J2	U29_J1	V+12	0.060706000000	0.049022000000
*J3	U29_J1	V+12	0.061976000000	0.049022000000
*K1	U29_J1	V+12	0.059436000000	0.047752000000
*K2	U29_J1	V+12	0.060706000000	0.047752000000
*K3	U29_J1	V+12	0.061976000000	0.047752000000
*L1	U29_J1	V+12	0.059436000000	0.046482000000
*L2	U29_J1	V+12	0.060706000000	0.046482000000
*L3	U29_J1	V+12	0.061976000000	0.046482000000
*L5	U29_J1	V+12	0.064516000000	0.046482000000
*[Ground Nets]
*A5	U29_L7	GND_DIGITAL	0.064516000000	0.059182000000
*A6	U29_L7	GND_DIGITAL	0.065786000000	0.059182000000
*A7	U29_L7	GND_DIGITAL	0.067056000000	0.059182000000
*B5	U29_L7	GND_DIGITAL	0.064516000000	0.057912000000
*B6	U29_L7	GND_DIGITAL	0.065786000000	0.057912000000
*B7	U29_L7	GND_DIGITAL	0.067056000000	0.057912000000
*C5	U29_L7	GND_DIGITAL	0.064516000000	0.056642000000
*C6	U29_L7	GND_DIGITAL	0.065786000000	0.056642000000
*C7	U29_L7	GND_DIGITAL	0.067056000000	0.056642000000
*D5	U29_L7	GND_DIGITAL	0.064516000000	0.055372000000
*D6	U29_L7	GND_DIGITAL	0.065786000000	0.055372000000
*D7	U29_L7	GND_DIGITAL	0.067056000000	0.055372000000
*E1	U29_L7	GND_DIGITAL	0.059436000000	0.054102000000
*E2	U29_L7	GND_DIGITAL	0.060706000000	0.054102000000
*E3	U29_L7	GND_DIGITAL	0.061976000000	0.054102000000
*E4	U29_L7	GND_DIGITAL	0.063246000000	0.054102000000
*E5	U29_L7	GND_DIGITAL	0.064516000000	0.054102000000
*E6	U29_L7	GND_DIGITAL	0.065786000000	0.054102000000
*E7	U29_L7	GND_DIGITAL	0.067056000000	0.054102000000
*F1	U29_L7	GND_DIGITAL	0.059436000000	0.052832000000
*F2	U29_L7	GND_DIGITAL	0.060706000000	0.052832000000
*F3	U29_L7	GND_DIGITAL	0.061976000000	0.052832000000
*F4	U29_L7	GND_DIGITAL	0.063246000000	0.052832000000
*F5	U29_L7	GND_DIGITAL	0.064516000000	0.052832000000
*F6	U29_L7	GND_DIGITAL	0.065786000000	0.052832000000
*F7	U29_L7	GND_DIGITAL	0.067056000000	0.052832000000
*G1	U29_L7	GND_DIGITAL	0.059436000000	0.051562000000
*G2	U29_L7	GND_DIGITAL	0.060706000000	0.051562000000
*G3	U29_L7	GND_DIGITAL	0.061976000000	0.051562000000
*G4	U29_L7	GND_DIGITAL	0.063246000000	0.051562000000
*G6	U29_L7	GND_DIGITAL	0.065786000000	0.051562000000
*H6	U29_L7	GND_DIGITAL	0.065786000000	0.050292000000
*J5	U29_L7	GND_DIGITAL	0.064516000000	0.049022000000
*J6	U29_L7	GND_DIGITAL	0.065786000000	0.049022000000
*K5	U29_L7	GND_DIGITAL	0.064516000000	0.047752000000
*K6	U29_L7	GND_DIGITAL	0.065786000000	0.047752000000
*L6	U29_L7	GND_DIGITAL	0.065786000000	0.046482000000
*L7	U29_L7	GND_DIGITAL	0.067056000000	0.046482000000
*
*
*[REM]***********************************************************************
*[Connection] U3 LM78L05_SO8_SOIC127P600X175-8N_IC_L78L08ACD13TR_PSL-00000009_L78L08ACD13TR 5
*[Connection Type] 
*[Power Nets]
*8	U3_8	V+12	0.004099000000	0.016518000000
*[Ground Nets]
*2	U3_3	GND_DIGITAL	0.009499000000	0.017788000000
*3	U3_3	GND_DIGITAL	0.009499000000	0.019058000000
*6	U3_3	GND_DIGITAL	0.004099000000	0.019058000000
*7	U3_3	GND_DIGITAL	0.004099000000	0.017788000000
*
*
*[REM]***********************************************************************
*[Connection] U30 LTM8025_LTUMODULE7X11_IC_LTM8025EV#PBF_PSL-00000026_LTM8025EV#PBF 65
*[Connection Type] 
*[Power Nets]
*A1	U30_A1	2V5	0.068834000000	0.059182000000
*A2	U30_A1	2V5	0.070104000000	0.059182000000
*A3	U30_A1	2V5	0.071374000000	0.059182000000
*A4	U30_A1	2V5	0.072644000000	0.059182000000
*B1	U30_A1	2V5	0.068834000000	0.057912000000
*B2	U30_A1	2V5	0.070104000000	0.057912000000
*B3	U30_A1	2V5	0.071374000000	0.057912000000
*B4	U30_A1	2V5	0.072644000000	0.057912000000
*C1	U30_A1	2V5	0.068834000000	0.056642000000
*C2	U30_A1	2V5	0.070104000000	0.056642000000
*C3	U30_A1	2V5	0.071374000000	0.056642000000
*C4	U30_A1	2V5	0.072644000000	0.056642000000
*D1	U30_A1	2V5	0.068834000000	0.055372000000
*D2	U30_A1	2V5	0.070104000000	0.055372000000
*D3	U30_A1	2V5	0.071374000000	0.055372000000
*D4	U30_A1	2V5	0.072644000000	0.055372000000
*H5	U30_H5	3V3	0.073914000000	0.050292000000
*J1	U30_J1	V+12	0.068834000000	0.049022000000
*J2	U30_J1	V+12	0.070104000000	0.049022000000
*J3	U30_J1	V+12	0.071374000000	0.049022000000
*K1	U30_J1	V+12	0.068834000000	0.047752000000
*K2	U30_J1	V+12	0.070104000000	0.047752000000
*K3	U30_J1	V+12	0.071374000000	0.047752000000
*L1	U30_J1	V+12	0.068834000000	0.046482000000
*L2	U30_J1	V+12	0.070104000000	0.046482000000
*L3	U30_J1	V+12	0.071374000000	0.046482000000
*L5	U30_J1	V+12	0.073914000000	0.046482000000
*[Ground Nets]
*A5	U30_A5	GND_DIGITAL	0.073914000000	0.059182000000
*A6	U30_A5	GND_DIGITAL	0.075184000000	0.059182000000
*A7	U30_A5	GND_DIGITAL	0.076454000000	0.059182000000
*B5	U30_A5	GND_DIGITAL	0.073914000000	0.057912000000
*B6	U30_A5	GND_DIGITAL	0.075184000000	0.057912000000
*B7	U30_A5	GND_DIGITAL	0.076454000000	0.057912000000
*C5	U30_A5	GND_DIGITAL	0.073914000000	0.056642000000
*C6	U30_A5	GND_DIGITAL	0.075184000000	0.056642000000
*C7	U30_A5	GND_DIGITAL	0.076454000000	0.056642000000
*D5	U30_A5	GND_DIGITAL	0.073914000000	0.055372000000
*D6	U30_A5	GND_DIGITAL	0.075184000000	0.055372000000
*D7	U30_A5	GND_DIGITAL	0.076454000000	0.055372000000
*E1	U30_A5	GND_DIGITAL	0.068834000000	0.054102000000
*E2	U30_A5	GND_DIGITAL	0.070104000000	0.054102000000
*E3	U30_A5	GND_DIGITAL	0.071374000000	0.054102000000
*E4	U30_A5	GND_DIGITAL	0.072644000000	0.054102000000
*E5	U30_A5	GND_DIGITAL	0.073914000000	0.054102000000
*E6	U30_A5	GND_DIGITAL	0.075184000000	0.054102000000
*E7	U30_A5	GND_DIGITAL	0.076454000000	0.054102000000
*F1	U30_A5	GND_DIGITAL	0.068834000000	0.052832000000
*F2	U30_A5	GND_DIGITAL	0.070104000000	0.052832000000
*F3	U30_A5	GND_DIGITAL	0.071374000000	0.052832000000
*F4	U30_A5	GND_DIGITAL	0.072644000000	0.052832000000
*F5	U30_A5	GND_DIGITAL	0.073914000000	0.052832000000
*F6	U30_A5	GND_DIGITAL	0.075184000000	0.052832000000
*F7	U30_A5	GND_DIGITAL	0.076454000000	0.052832000000
*G1	U30_A5	GND_DIGITAL	0.068834000000	0.051562000000
*G2	U30_A5	GND_DIGITAL	0.070104000000	0.051562000000
*G3	U30_A5	GND_DIGITAL	0.071374000000	0.051562000000
*G4	U30_A5	GND_DIGITAL	0.072644000000	0.051562000000
*G6	U30_A5	GND_DIGITAL	0.075184000000	0.051562000000
*H6	U30_A5	GND_DIGITAL	0.075184000000	0.050292000000
*J5	U30_A5	GND_DIGITAL	0.073914000000	0.049022000000
*J6	U30_A5	GND_DIGITAL	0.075184000000	0.049022000000
*K5	U30_A5	GND_DIGITAL	0.073914000000	0.047752000000
*K6	U30_A5	GND_DIGITAL	0.075184000000	0.047752000000
*L6	U30_A5	GND_DIGITAL	0.075184000000	0.046482000000
*L7	U30_A5	GND_DIGITAL	0.076454000000	0.046482000000
*
*
*[REM]***********************************************************************
*[Connection] U31 LTM8025_LTUMODULE7X11_IC_LTM8025EV#PBF_PSL-00000026_LTM8025EV#PBF 64
*[Connection Type] 
*[Power Nets]
*A1	U31_A1	3V3	0.078232000000	0.059182000000
*A2	U31_A1	3V3	0.079502000000	0.059182000000
*A3	U31_A1	3V3	0.080772000000	0.059182000000
*A4	U31_A1	3V3	0.082042000000	0.059182000000
*B1	U31_A1	3V3	0.078232000000	0.057912000000
*B2	U31_A1	3V3	0.079502000000	0.057912000000
*B3	U31_A1	3V3	0.080772000000	0.057912000000
*B4	U31_A1	3V3	0.082042000000	0.057912000000
*C1	U31_A1	3V3	0.078232000000	0.056642000000
*C2	U31_A1	3V3	0.079502000000	0.056642000000
*C3	U31_A1	3V3	0.080772000000	0.056642000000
*C4	U31_A1	3V3	0.082042000000	0.056642000000
*D1	U31_A1	3V3	0.078232000000	0.055372000000
*D2	U31_A1	3V3	0.079502000000	0.055372000000
*D3	U31_A1	3V3	0.080772000000	0.055372000000
*D4	U31_A1	3V3	0.082042000000	0.055372000000
*J1	U31_J1	V+12	0.078232000000	0.049022000000
*J2	U31_J1	V+12	0.079502000000	0.049022000000
*J3	U31_J1	V+12	0.080772000000	0.049022000000
*K1	U31_J1	V+12	0.078232000000	0.047752000000
*K2	U31_J1	V+12	0.079502000000	0.047752000000
*K3	U31_J1	V+12	0.080772000000	0.047752000000
*L1	U31_J1	V+12	0.078232000000	0.046482000000
*L2	U31_J1	V+12	0.079502000000	0.046482000000
*L3	U31_J1	V+12	0.080772000000	0.046482000000
*L5	U31_J1	V+12	0.083312000000	0.046482000000
*[Ground Nets]
*A5	U31_L7	GND_DIGITAL	0.083312000000	0.059182000000
*A6	U31_L7	GND_DIGITAL	0.084582000000	0.059182000000
*A7	U31_L7	GND_DIGITAL	0.085852000000	0.059182000000
*B5	U31_L7	GND_DIGITAL	0.083312000000	0.057912000000
*B6	U31_L7	GND_DIGITAL	0.084582000000	0.057912000000
*B7	U31_L7	GND_DIGITAL	0.085852000000	0.057912000000
*C5	U31_L7	GND_DIGITAL	0.083312000000	0.056642000000
*C6	U31_L7	GND_DIGITAL	0.084582000000	0.056642000000
*C7	U31_L7	GND_DIGITAL	0.085852000000	0.056642000000
*D5	U31_L7	GND_DIGITAL	0.083312000000	0.055372000000
*D6	U31_L7	GND_DIGITAL	0.084582000000	0.055372000000
*D7	U31_L7	GND_DIGITAL	0.085852000000	0.055372000000
*E1	U31_L7	GND_DIGITAL	0.078232000000	0.054102000000
*E2	U31_L7	GND_DIGITAL	0.079502000000	0.054102000000
*E3	U31_L7	GND_DIGITAL	0.080772000000	0.054102000000
*E4	U31_L7	GND_DIGITAL	0.082042000000	0.054102000000
*E5	U31_L7	GND_DIGITAL	0.083312000000	0.054102000000
*E6	U31_L7	GND_DIGITAL	0.084582000000	0.054102000000
*E7	U31_L7	GND_DIGITAL	0.085852000000	0.054102000000
*F1	U31_L7	GND_DIGITAL	0.078232000000	0.052832000000
*F2	U31_L7	GND_DIGITAL	0.079502000000	0.052832000000
*F3	U31_L7	GND_DIGITAL	0.080772000000	0.052832000000
*F4	U31_L7	GND_DIGITAL	0.082042000000	0.052832000000
*F5	U31_L7	GND_DIGITAL	0.083312000000	0.052832000000
*F6	U31_L7	GND_DIGITAL	0.084582000000	0.052832000000
*F7	U31_L7	GND_DIGITAL	0.085852000000	0.052832000000
*G1	U31_L7	GND_DIGITAL	0.078232000000	0.051562000000
*G2	U31_L7	GND_DIGITAL	0.079502000000	0.051562000000
*G3	U31_L7	GND_DIGITAL	0.080772000000	0.051562000000
*G4	U31_L7	GND_DIGITAL	0.082042000000	0.051562000000
*G6	U31_L7	GND_DIGITAL	0.084582000000	0.051562000000
*H6	U31_L7	GND_DIGITAL	0.084582000000	0.050292000000
*J5	U31_L7	GND_DIGITAL	0.083312000000	0.049022000000
*J6	U31_L7	GND_DIGITAL	0.084582000000	0.049022000000
*K5	U31_L7	GND_DIGITAL	0.083312000000	0.047752000000
*K6	U31_L7	GND_DIGITAL	0.084582000000	0.047752000000
*L6	U31_L7	GND_DIGITAL	0.084582000000	0.046482000000
*L7	U31_L7	GND_DIGITAL	0.085852000000	0.046482000000
*
*
*[REM]***********************************************************************
*[Connection] U32 TLC5602A_SOIC127P1028X265-20N_IC_TLC5602CDWR_PSL-00000028_TLC5602CDWR 7
*[Connection Type] 
*[Power Nets]
*2	U32_2	VCC	0.066731000000	-0.001348000000
*9	U32_2	VCC	0.066731000000	0.007542000000
*[Ground Nets]
*1	U32_10	GND_DIGITAL	0.066731000000	-0.002618000000
*10	U32_10	GND_DIGITAL	0.066731000000	0.008812000000
*20	U32_10	GND_DIGITAL	0.057331000000	-0.002618000000
*3	U32_10	GND_DIGITAL	0.066731000000	-0.000078000000
*7	U32_10	GND_DIGITAL	0.066731000000	0.005002000000
*
*
*[REM]***********************************************************************
*[Connection] U33 DG419A_SOG0508WG244L225_IC_DG419CY+_PSL-00000008_DG419CY+ 3
*[Connection Type] 
*[Power Nets]
*4	U33_4	V+12	0.075031000000	0.008507000000
*7	U33_7	V12N	0.070053000000	0.005967000000
*[Ground Nets]
*3	U33_3	GND_DIGITAL	0.075031000000	0.007237000000
*
*[REM]***********************************************************************
*[Connection] U35 TLC5602A_SOIC127P1028X265-20N_IC_TLC5602CDWR_PSL-00000028_TLC5602CDWR 7
*[Connection Type] 
*[Power Nets]
*2	U35_9	VCC	0.066731000000	0.014130000000
*9	U35_9	VCC	0.066731000000	0.023020000000
*[Ground Nets]
*1	U35_10	GND_DIGITAL	0.066731000000	0.012860000000
*10	U35_10	GND_DIGITAL	0.066731000000	0.024290000000
*20	U35_10	GND_DIGITAL	0.057331000000	0.012860000000
*3	U35_10	GND_DIGITAL	0.066731000000	0.015400000000
*7	U35_10	GND_DIGITAL	0.066731000000	0.020480000000
*
*
*[REM]***********************************************************************
*[Connection] U36 DG419A_SOG0508WG244L225_IC_DG419CY+_PSL-00000008_DG419CY+ 3
*[Connection Type] 
*[Power Nets]
*4	U36_4	V+12	0.075031000000	0.023985000000
*7	U36_7	V12N	0.070053000000	0.021445000000
*[Ground Nets]
*3	U36_3	GND_DIGITAL	0.075031000000	0.022715000000
*
*[REM]***********************************************************************
*[Connection] U38 FF_D_8X_OE3S_20P_SOIC127P1032X265-20AN_IC_74HCT574_EMA-00007307V22_74HCT574 3
*[Connection Type] 
*[Power Nets]
*20	U38_20	VCC	0.053195000000	0.008814000000
*[Ground Nets]
*1	U38_1	GND_DIGITAL	0.043695000000	0.008814000000
*10	U38_1	GND_DIGITAL	0.043695000000	-0.002616000000
*
*
*[REM]***********************************************************************
*[Connection] U39 FF_D_8X_OE3S_20P_SOIC127P1032X265-20AN_IC_74HCT574_EMA-00007307V22_74HCT574 3
*[Connection Type] 
*[Power Nets]
*20	U39_20	VCC	0.053195000000	0.024292000000
*[Ground Nets]
*1	U39_1	GND_DIGITAL	0.043695000000	0.024292000000
*10	U39_1	GND_DIGITAL	0.043695000000	0.012862000000
*
*
*[REM]***********************************************************************
*[Connection] U40 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U40_32	VCC	0.012813000000	0.109220000000
*[Ground Nets]
*16	U40_16	GND_DIGITAL	0.005713000000	0.090170000000
*24	U40_16	GND_DIGITAL	0.012813000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U41 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U41_32	VCC	0.023727000000	0.109220000000
*[Ground Nets]
*16	U41_16	GND_DIGITAL	0.016627000000	0.090170000000
*24	U41_16	GND_DIGITAL	0.023727000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U42 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U42_32	VCC	0.034641000000	0.109220000000
*[Ground Nets]
*16	U42_24	GND_DIGITAL	0.027541000000	0.090170000000
*24	U42_24	GND_DIGITAL	0.034641000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U43 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U43_32	VCC	0.045555000000	0.109220000000
*[Ground Nets]
*16	U43_24	GND_DIGITAL	0.038455000000	0.090170000000
*24	U43_24	GND_DIGITAL	0.045555000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U44 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U44_32	VCC	0.056469000000	0.109220000000
*[Ground Nets]
*16	U44_24	GND_DIGITAL	0.049369000000	0.090170000000
*24	U44_24	GND_DIGITAL	0.056469000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U45 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U45_32	VCC	0.067383000000	0.109220000000
*[Ground Nets]
*16	U45_16	GND_DIGITAL	0.060283000000	0.090170000000
*24	U45_16	GND_DIGITAL	0.067383000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U46 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U46_32	VCC	0.078297000000	0.109220000000
*[Ground Nets]
*16	U46_16	GND_DIGITAL	0.071197000000	0.090170000000
*24	U46_16	GND_DIGITAL	0.078297000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U47 UPD431000AGW-B15_SOJ127P866X375-32N_IC_UPD431000AGW-B15_PSL-00000035_UPD431000AGW-B15 3
*[Connection Type] 
*[Power Nets]
*32	U47_32	VCC	0.089211000000	0.109220000000
*[Ground Nets]
*16	U47_16	GND_DIGITAL	0.082111000000	0.090170000000
*24	U47_16	GND_DIGITAL	0.089211000000	0.099060000000
*
*
*[REM]***********************************************************************
*[Connection] U48 74-245_20P_SOIC127P1028X265-20N_IC_74ACT245_EMA-00006591V22_74ACT245 2
*[Connection Type] 
*[Power Nets]
*20	U48_20	VCC	0.000636000000	0.019939000000
*[Ground Nets]
*10	U48_10	GND_DIGITAL	-0.008764000000	0.008509000000
*
*[REM]***********************************************************************
*[Connection] U49 MAX6711_SOT343N_IC_MAX6711S_EMA-00006895V22_MAX6711S 2
*[Connection Type] 
*[Power Nets]
*4	U49_4	VCC	0.040016000000	0.025415000000
*[Ground Nets]
*1	U49_1	GND_DIGITAL	0.038216000000	0.025415000000
*
*[REM]***********************************************************************
*[Connection] U5 VREG_TGND_TO254P1410X464-4N_IC_LM340_EMA-00007000V22_LM340 3
*[Connection Type] 
*[Power Nets]
*1	U5_1	V+12	0.012106000000	0.011523000000
*[Ground Nets]
*2	U5_4	GND_DIGITAL	0.009566000000	0.011523000000
*4	U5_4	GND_DIGITAL	0.009566000000	0.001423000000
*
*
*[REM]***********************************************************************
*[Connection] U50 NBC12429_QFN50P500X500X100-33N_IC_NBC12429AMNR4G_PSL-00000017_NBC12429AMNR4G 18
*[Connection Type] 
*[Power Nets]
*27	U50_28	VCC	0.042480000000	0.029095000000
*28	U50_28	VCC	0.042480000000	0.029595000000
*32	U50_28	VCC	0.042480000000	0.031595000000
*[Ground Nets]
*1	U50_1	GND_DIGITAL	0.041755000000	0.032320000000
*12	U50_1	GND_DIGITAL	0.037530000000	0.030095000000
*13	U50_1	GND_DIGITAL	0.037530000000	0.029595000000
*14	U50_1	GND_DIGITAL	0.037530000000	0.029095000000
*15	U50_1	GND_DIGITAL	0.037530000000	0.028595000000
*17	U50_1	GND_DIGITAL	0.038255000000	0.027370000000
*18	U50_1	GND_DIGITAL	0.038755000000	0.027370000000
*2	U50_1	GND_DIGITAL	0.041255000000	0.032320000000
*20	U50_1	GND_DIGITAL	0.039755000000	0.027370000000
*22	U50_1	GND_DIGITAL	0.040755000000	0.027370000000
*23	U50_1	GND_DIGITAL	0.041255000000	0.027370000000
*25	U50_1	GND_DIGITAL	0.042480000000	0.028095000000
*29	U50_1	GND_DIGITAL	0.042480000000	0.030095000000
*3	U50_1	GND_DIGITAL	0.040755000000	0.032320000000
*33	U50_1	GND_DIGITAL	0.040005000000	0.029845000000
*
*
*[REM]***********************************************************************
*[Connection] U51 TPS51200_DRC10_2P4X1P65_IC_TPS51200DRCR_PSL-00000036_TPS51200DRCR 7
*[Connection Type] 
*[Power Nets]
*10	U51_10	3V3	0.048719000000	0.031099000000
*7	U51_10	3V3	0.048719000000	0.029599000000
*2	U51_2	1V8	0.045769000000	0.030599000000
*3	U51_5	0V9	0.045769000000	0.030099000000
*5	U51_5	0V9	0.045769000000	0.029099000000
*[Ground Nets]
*4	U51_8	GND_DIGITAL	0.045769000000	0.029599000000
*8	U51_8	GND_DIGITAL	0.048719000000	0.030099000000
*
*
*[REM]***********************************************************************
*[Connection] U6 FCT16245_SOP50P810X110-48N_IC_74ALVT16245DGG_118_PSL-00000016_0_0_0_0_74ALVT16245DGG_118 14
*[Connection Type] 
*[Power Nets]
*18	U6_42	VCC	-0.007356000000	0.078657000000
*31	U6_42	VCC	0.000244000000	0.078657000000
*42	U6_42	VCC	0.000244000000	0.084157000000
*7	U6_42	VCC	-0.007356000000	0.084157000000
*[Ground Nets]
*10	U6_25	GND_DIGITAL	-0.007356000000	0.082657000000
*15	U6_25	GND_DIGITAL	-0.007356000000	0.080157000000
*21	U6_25	GND_DIGITAL	-0.007356000000	0.077157000000
*24	U6_25	GND_DIGITAL	-0.007356000000	0.075657000000
*25	U6_25	GND_DIGITAL	0.000244000000	0.075657000000
*28	U6_25	GND_DIGITAL	0.000244000000	0.077157000000
*34	U6_25	GND_DIGITAL	0.000244000000	0.080157000000
*39	U6_25	GND_DIGITAL	0.000244000000	0.082657000000
*4	U6_25	GND_DIGITAL	-0.007356000000	0.085657000000
*45	U6_25	GND_DIGITAL	0.000244000000	0.085657000000
*
*
*[REM]***********************************************************************
*[Connection] U7 74-245_20P_SOIC127P1028X265-20N_IC_74ACT245_EMA-00006591V22_74ACT245 2
*[Connection Type] 
*[Power Nets]
*20	U7_20	VCC	0.000636000000	0.035179000000
*[Ground Nets]
*10	U7_10	GND_DIGITAL	-0.008764000000	0.023749000000
*
*[REM]***********************************************************************
*[Connection] U8 FCT16245_SOP50P810X110-48N_IC_74ALVT16245DGG_118_PSL-00000016_0_0_0_0_74ALVT16245DGG_118 14
*[Connection Type] 
*[Power Nets]
*18	U8_42	VCC	-0.007356000000	0.061893000000
*31	U8_42	VCC	0.000244000000	0.061893000000
*42	U8_42	VCC	0.000244000000	0.067393000000
*7	U8_42	VCC	-0.007356000000	0.067393000000
*[Ground Nets]
*1	U8_34	GND_DIGITAL	-0.007356000000	0.070393000000
*10	U8_34	GND_DIGITAL	-0.007356000000	0.065893000000
*15	U8_34	GND_DIGITAL	-0.007356000000	0.063393000000
*21	U8_34	GND_DIGITAL	-0.007356000000	0.060393000000
*28	U8_34	GND_DIGITAL	0.000244000000	0.060393000000
*34	U8_34	GND_DIGITAL	0.000244000000	0.063393000000
*39	U8_34	GND_DIGITAL	0.000244000000	0.065893000000
*4	U8_34	GND_DIGITAL	-0.007356000000	0.068893000000
*45	U8_34	GND_DIGITAL	0.000244000000	0.068893000000
*48	U8_34	GND_DIGITAL	0.000244000000	0.070393000000
*
*
*[REM]***********************************************************************
*[Connection] U9 FCT16245_SOP50P810X110-48N_IC_74ALVT16245DGG_118_PSL-00000016_0_0_0_0_74ALVT16245DGG_118 14
*[Connection Type] 
*[Power Nets]
*18	U9_42	VCC	-0.007483000000	0.044875000000
*31	U9_42	VCC	0.000117000000	0.044875000000
*42	U9_42	VCC	0.000117000000	0.050375000000
*7	U9_42	VCC	-0.007483000000	0.050375000000
*[Ground Nets]
*10	U9_4	GND_DIGITAL	-0.007483000000	0.048875000000
*15	U9_4	GND_DIGITAL	-0.007483000000	0.046375000000
*21	U9_4	GND_DIGITAL	-0.007483000000	0.043375000000
*24	U9_4	GND_DIGITAL	-0.007483000000	0.041875000000
*25	U9_4	GND_DIGITAL	0.000117000000	0.041875000000
*28	U9_4	GND_DIGITAL	0.000117000000	0.043375000000
*34	U9_4	GND_DIGITAL	0.000117000000	0.046375000000
*39	U9_4	GND_DIGITAL	0.000117000000	0.048875000000
*4	U9_4	GND_DIGITAL	-0.007483000000	0.051875000000
*45	U9_4	GND_DIGITAL	0.000117000000	0.051875000000
*
*
*[REM]***********************************************************************
*[Connection] zakorotka_01 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	J6_A1	V+12	-0.012784000000	0.025285000000
*[Ground Nets]
*2	J6_C1	GND_DIGITAL	-0.016284000000	0.025795000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_02 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	J6_D3	V12N	-0.012784000000	0.028335000000
*[Ground Nets]
*2	J6_C1	GND_DIGITAL	-0.016284000000	0.027825000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_03 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*2	P1_2	0V9	0.024900000000	0.025860000000
*[Ground Nets]
*1	P1_1	GND_DIGITAL	0.024900000000	0.028400000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_04 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*2	P1_4	1V2	0.022360000000	0.025860000000
*[Ground Nets]
*1	P1_1	GND_DIGITAL	0.019820000000	0.028400000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_05 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	P1_6	1V8	0.019820000000	0.025860000000
*[Ground Nets]
*2	P1_1	GND_DIGITAL	0.019820000000	0.028400000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_06 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	P1_14	2V5	0.009660000000	0.025860000000
*[Ground Nets]
*2	P1_1	GND_DIGITAL	0.009660000000	0.028400000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_07 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*2	U29_J1	V+12	0.061976000000	0.049022000000
*[Ground Nets]
*1	U29_L7	GND_DIGITAL	0.064516000000	0.049022000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_08 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	U29_H5	3V3	0.064516000000	0.050292000000
*[Ground Nets]
*2	U29_L7	GND_DIGITAL	0.065786000000	0.050292000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_09 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	U30_A1	2V5	0.072644000000	0.055372000000
*[Ground Nets]
*2	U30_A5	GND_DIGITAL	0.073914000000	0.055372000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_10 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	U31_J1	V+12	0.080772000000	0.049022000000
*[Ground Nets]
*2	U31_L7	GND_DIGITAL	0.083312000000	0.049022000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_11 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	U31_A1	3V3	0.082042000000	0.055372000000
*[Ground Nets]
*2	U31_L7	GND_DIGITAL	0.083312000000	0.055372000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_12 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	U30_H5	3V3	0.073914000000	0.050292000000
*[Ground Nets]
*2	U30_A5	GND_DIGITAL	0.075184000000	0.050292000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_13 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	U30_J1	V+12	0.073914000000	0.046482000000
*[Ground Nets]
*2	U30_A5	GND_DIGITAL	0.073914000000	0.047752000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_14 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	U29_A1	1V2	0.063246000000	0.055372000000
*[Ground Nets]
*2	U29_L7	GND_DIGITAL	0.064516000000	0.055372000000
*
*[REM]***********************************************************************
*[Connection] zakorotka_15 Zakorotka 2
*[Connection Type] 
*[Power Nets]
*1	J6_A23	VCC	-0.012784000000	0.079135000000
*[Ground Nets]
*2	J6_C1	GND_DIGITAL	-0.016284000000	0.081675000000
*
*[MCP End]
*
*This concludes the MCP section
*Define the S element, the Model file is output from BNP

.MODEL   Spara   S		
+		BNPFILE = "Cadence_Demo_091724_163748_8672.BNP"

S		
+			J5_1	J5_4
+			J6_A1	J6_C1
+			J6_D3	J6_C1
+			J6_A23	J6_C1
+			J7_137	J7_99
+			LCD1_2	LCD1_1
+			LCD2_2	LCD2_1
+			P1_2	P1_1
+			P1_4	P1_1
+			P1_6	P1_1
+			P1_14	P1_1
+			P1_12	P1_1
+			U1_K10	U1_T1
+			U1_R4	U1_T1
+			U1_D15	U1_T1
+			U2_K10	U2_A16
+			U2_B13	U2_A16
+			U2_R8	U2_A16
+			U2_K13	U2_A16
+			U3_8	U3_3
+			U5_1	U5_4
+			U6_42	U6_25
+			U7_20	U7_10
+			U8_42	U8_34
+			U9_42	U9_4
+			U10_20	U10_11
+			U10_18	U10_11
+			U11_20	U11_11
+			U11_18	U11_11
+			U12_J2	U12_N1
+			U12_A9	U12_N1
+			U13_J2	U13_B2
+			U13_A1	U13_B2
+			U22_20	U22_1
+			U29_A1	U29_L7
+			U29_H5	U29_L7
+			U29_J1	U29_L7
+			U30_A1	U30_A5
+			U30_H5	U30_A5
+			U30_J1	U30_A5
+			U31_A1	U31_L7
+			U31_J1	U31_L7
+			U32_2	U32_10
+			U33_4	U33_3
+			U33_7	U33_3
+			U35_9	U35_10
+			U36_4	U36_3
+			U36_7	U36_3
+			U38_20	U38_1
+			U39_20	U39_1
+			U40_32	U40_16
+			U41_32	U41_16
+			U42_32	U42_24
+			U43_32	U43_24
+			U44_32	U44_24
+			U45_32	U45_16
+			U46_32	U46_16
+			U47_32	U47_16
+			U48_20	U48_10
+			U49_4	U49_1
+			U50_28	U50_1
+			U51_5	U51_8
+			U51_2	U51_8
+			U51_10	U51_8
+			MNAME = Spara

*
.ENDS
*